module datapath(
	// Port Declarations
);

	// File for Creating the Datapath

endmodule
