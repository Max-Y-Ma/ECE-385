module ripple_adder_4bit (
	input  [3:0] A, B,
	input         cin,
	output [3:0] S,
	output        cout
);

    /* TODO
     *
     * Insert code here to implement a 4 bit ripple adder.
	  * To be used for 16 bit ripple adder and carry-select adder
     * Your code should be completly combinational (don't use always_ff or always_latch).
     * Feel free to create sub-modules or other files. */

     
endmodule