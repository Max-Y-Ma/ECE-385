//control_unit (
//
//	);
//
//endmodule
